library ieee;
use ieee.std_logic_1164.all;

entity sub_4bit is
  port(
    A, B  : in  std_logic_vector(3 downto 0);
    Bin   : in  std_logic;                     -- De forma inicial 0
    D     : out std_logic_vector(3 downto 0);  -- diferencia
    Bout  : out std_logic                      -- prestamos en casos que se salga
  );
end entity;

architecture structural of sub_4bit is			-- Structural para unir componenetes mas pequeños
  component full_sub_1bit
    port(A,B,Bin: in std_logic; D,Bout: out std_logic);	-- Entradas y salidas
  end component;

  signal b1,b2,b3: std_logic;  -- Prestamo internos
begin
  u0: full_sub_1bit port map(A=>A(0), B=>B(0), Bin=>Bin, D=>D(0), Bout=>b1);
  u1: full_sub_1bit port map(A=>A(1), B=>B(1), Bin=>b1 , D=>D(1), Bout=>b2);
  u2: full_sub_1bit port map(A=>A(2), B=>B(2), Bin=>b2 , D=>D(2), Bout=>b3);
  u3: full_sub_1bit port map(A=>A(3), B=>B(3), Bin=>b3 , D=>D(3), Bout=>Bout);
end architecture;
